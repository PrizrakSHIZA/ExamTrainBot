    ����          CExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null   �System.Collections.Generic.List`1[[ExamTrainBot.Tests.Test, ExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  ExamTrainBot.Tests.Test[]   	                   ExamTrainBot.Tests.Test   	   	      ExamTrainBot.Tests.Test   Text	questions�System.Collections.Generic.List`1[[ExamTrainBot.Tests.Questions.Question, ExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]      New test	            новый тест		      �System.Collections.Generic.List`1[[ExamTrainBot.Tests.Questions.Question, ExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  'ExamTrainBot.Tests.Questions.Question[]   	
         	      	         
          %ExamTrainBot.Tests.Questions.Question   	   	   	   
          %ExamTrainBot.Tests.Questions.Question   	      /ExamTrainBot.Tests.Questions.ConformityQuestion   <text>k__BackingField<points>k__BackingField<answer>k__BackingField<variants>k__BackingFieldruledelimiterChars       H1) 1
2) 2
3) 3
4) 4

А) один
Б) два
В) три
Г) чотири      1а 2б 3в 4г
   g
(Будь ласка заповнюйте відповідь у вигляді: 'А-1,Б-2,В-3,Г-4')	      )ExamTrainBot.Tests.Questions.TestQuestion   <text>k__BackingField<points>k__BackingField<variants>k__BackingFieldcolumns<answer>k__BackingField        ?   	         !   )ExamTrainBot.Tests.Questions.FreeQuestion   <text>k__BackingField<points>k__BackingField<answer>k__BackingField<variants>k__BackingFieldrule       Ви людина?      Так
   _
(Будь ласка, будьте уважні при написанні відповіді!)         Проверка   	         два       ,.	
         !   !!   ?    ??      !   один"   два#   три$   четыре