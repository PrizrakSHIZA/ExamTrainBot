    ����          CExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null   �System.Collections.Generic.List`1[[ExamTrainBot.Tests.Test, ExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  ExamTrainBot.Tests.Test[]   	                   ExamTrainBot.Tests.Test   	      ExamTrainBot.Tests.Test   Text	questions�System.Collections.Generic.List`1[[ExamTrainBot.Tests.Questions.Question, ExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]      Якесь правило.	      �System.Collections.Generic.List`1[[ExamTrainBot.Tests.Questions.Question, ExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  'ExamTrainBot.Tests.Questions.Question[]   	                   %ExamTrainBot.Tests.Questions.Question   	   		   	
   
   )ExamTrainBot.Tests.Questions.TestQuestion   <text>k__BackingField<points>k__BackingField<variants>k__BackingFieldcolumns<answer>k__BackingField        ?Питання 1 (Правильна відповідь це 2)    	         2	   )ExamTrainBot.Tests.Questions.FreeQuestion   <text>k__BackingField<points>k__BackingField<answer>k__BackingField<variants>k__BackingFieldrule       EПитання 2, вільне відповідь. Ви людина?       Так
   _
(Будь ласка, будьте уважні при написанні відповіді!)
   /ExamTrainBot.Tests.Questions.ConformityQuestion   <text>k__BackingField<points>k__BackingField<answer>k__BackingField<variants>k__BackingFieldruledelimiterChars       ~Питання 3(відповідність)
1) 1
2) 2
3) 3
4) 4

А) Один
Б) Два
В) Три
Г) Чотири       1а,б2,3в,г4
   g
(Будь ласка заповнюйте відповідь у вигляді: 'А-1,Б-2,В-3,Г-4')	            1   2   3   4       ,.	
