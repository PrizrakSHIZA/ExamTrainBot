    ����          CExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null   {System.Collections.Generic.List`1[[ExamTrainBot.User, ExamTrainBot, Version=1.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  ExamTrainBot.User[]   	                   ExamTrainBot.User   	      ExamTrainBot.User   idname
subscriberisadminontestpointscurrentquestiontestcreation       	   ��8=       Ефим Ряскин           